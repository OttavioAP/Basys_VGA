//top



